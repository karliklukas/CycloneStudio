module cLED0(input wire IN, output wire LED0);
//hidden: LED0
//position: 303,85,DE0nano
assign LED0 = IN;
endmodule
