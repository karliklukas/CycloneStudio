module cOUT_PIN10(input wire OUT, output wire PIN10);
//hidden: PIN10
assign PIN10 = OUT;
endmodule
