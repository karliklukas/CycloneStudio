module cTTre(input wire OUT, output wire TTre);
//hidden: TTre
assign TTre = OUT;
endmodule
