module cOUT_PIN9(input wire OUT, output wire PIN9);
//hidden: PIN9
assign PIN9 = OUT;
endmodule
