module cIN_PIN12(input wire IN_PIN12, output wire IN);
//hidden: IN_PIN12
assign IN = IN_PIN12;
endmodule
