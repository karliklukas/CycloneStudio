module cOUT_PIN1(input wire OUT, output wire OUT_PIN1);
//hidden: OUT_PIN1
//position: 129,37,DE0nano;195,396,StormIV
assign OUT_PIN1 = OUT;
endmodule
