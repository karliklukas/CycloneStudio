module cOUT_PIN2(input wire OUT, output wire OUT_PIN2);
//hidden: OUT_PIN2
//position: 143,37,DE0nano;195,407,StormIV
assign OUT_PIN2 = OUT;
endmodule
