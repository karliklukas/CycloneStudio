module cvystup5(input wire OUT, output wire vystup5);
//hidden: vystup5
assign vystup5 = OUT;
endmodule
