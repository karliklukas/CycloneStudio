module cIN_PIN16(input wire IN_PIN16, output wire IN);
//hidden: IN_PIN16
assign IN = IN_PIN16;
endmodule
