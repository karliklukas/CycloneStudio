module cIN_PIN4(input wire IN_PIN4, output wire IN);
//hidden: IN_PIN4
assign IN = IN_PIN4;
endmodule
