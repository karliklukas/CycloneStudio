module cOUT_PIN7(input wire OUT, output wire OUT_PIN7);
//hidden: OUT_PIN7
assign OUT_PIN7 = OUT;
endmodule
