module cOUT_PIN17(input wire OUT, output wire OUT_PIN17);
//hidden: OUT_PIN17
//position: 389,37,DE0nano
assign OUT_PIN17 = OUT;
endmodule
