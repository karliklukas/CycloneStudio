module cOUT_PIN17(input wire OUT, output wire OUT_PIN17);
//hidden: OUT_PIN17
assign OUT_PIN17 = OUT;
endmodule
