module cLED2(input wire IN, output wire LED2);
//hidden: LED2
//position: 110,368,StormIV
assign LED2 = IN;
endmodule
