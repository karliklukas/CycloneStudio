module cIN_PIN13(input wire IN_PIN13, output wire IN);
//hidden: IN_PIN13
//position: 317,300,DE0nano
assign IN = IN_PIN13;
endmodule
