module cOUT_PIN14(input wire OUT, output wire OUT_PIN14);
//hidden: OUT_PIN14
assign OUT_PIN14 = OUT;
endmodule
