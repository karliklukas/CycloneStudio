module cOUT_PIN19(input wire OUT, output wire OUT_PIN19);
//hidden: OUT_PIN19
assign OUT_PIN19 = OUT;
endmodule
