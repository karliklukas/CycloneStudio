module cLED8(input wire IN, output wire LED8);
//hidden: LED8
assign LED8 = IN;
endmodule
