module cOUT_PIN5(input wire OUT, output wire OUT_PIN5);
//hidden: OUT_PIN5
assign OUT_PIN5 = OUT;
endmodule
