module cLED6(input wire IN, output wire LED6);
//hidden: LED6
//position: 110,278,StormIV
assign LED6 = IN;
endmodule
