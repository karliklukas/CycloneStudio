module cinCLK(input wire inCLK, output wire IN);
//hidden: inCLK
assign IN = inCLK;
endmodule
