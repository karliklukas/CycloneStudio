module cOUT_PIN1(input wire OUT, output wire OUT_PIN1);
//hidden: OUT_PIN1
assign OUT_PIN1 = OUT;
endmodule
