module cLED4(input wire IN, output wire LED4);
//hidden: LED4
//position: 235,85,DE0nano
assign LED4 = IN;
endmodule
