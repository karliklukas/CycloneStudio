module cIN_PIN6(input wire IN_PIN6, output wire IN);
//hidden: IN_PIN6
//position: 216,300,DE0nano;281,196,StormIV
assign IN = IN_PIN6;
endmodule
