module cIN_PIN5(input wire PIN5, output wire IN);
//hidden: PIN5
assign IN = PIN5;
endmodule
