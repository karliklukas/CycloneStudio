module cIN_PIN19(input wire IN_PIN19, output wire IN);
//hidden: IN_PIN19
assign IN = IN_PIN19;
endmodule
