module cOUT_PIN6(input wire OUT, output wire PIN6);
//hidden: PIN6
assign PIN6 = OUT;
endmodule
