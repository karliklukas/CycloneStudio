module cONE(output wire Y);
assign Y = 1'b1;
endmodule
