module cOUT_PIN8(input wire OUT, output wire OUT_PIN8);
//hidden: OUT_PIN8
//position: 244,37,DE0nano;227,407,StormIV
assign OUT_PIN8 = OUT;
endmodule
