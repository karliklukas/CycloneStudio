module cKEY0(input wire KEY0, output wire OUT);
//hidden: KEY0
assign OUT = KEY0;
endmodule
