module cOUT_PIN20(input wire OUT, output wire OUT_PIN20);
//hidden: OUT_PIN20
//position: 389,51,DE0nano
assign OUT_PIN20 = OUT;
endmodule
