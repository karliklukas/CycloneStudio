module cIN_PIN3(input wire IN_PIN3, output wire IN);
//hidden: IN_PIN3
assign IN = IN_PIN3;
endmodule
