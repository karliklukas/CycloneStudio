module cIN_PIN2(input wire PIN2, output wire IN);
//hidden: PIN2
assign IN = PIN2;
endmodule
