module cKEY3(input wire KEY3, output wire OUT);
//hidden: KEY3
assign OUT = KEY3;
endmodule
