module cvstup1(input wire vstup1, output wire IN);
//hidden: vstup1
assign IN = vstup1;
endmodule
