module cLED6(input wire IN, output wire LED6);
//hidden: LED6
assign LED6 = IN;
endmodule
