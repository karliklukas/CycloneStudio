module cIN_PIN17(input wire IN_PIN17, output wire IN);
//hidden: IN_PIN17
assign IN = IN_PIN17;
endmodule
