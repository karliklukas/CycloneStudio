module cout_LED0(input wire OUT, output wire out_LED0);
//hidden: out_LED0
assign out_LED0 = OUT;
endmodule
