module cCustOut(input wire OUT, output wire CustOut);
//hidden: CustOut
assign CustOut = OUT;
endmodule
