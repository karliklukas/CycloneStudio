module cvstup2(input wire vstup2, output wire IN);
//hidden: vstup2
assign IN = vstup2;
endmodule
