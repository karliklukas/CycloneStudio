module cvystup1(input wire OUT, output wire vystup1);
//hidden: vystup1
assign vystup1 = OUT;
endmodule
