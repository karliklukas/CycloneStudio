module cLED5(input wire IN, output wire LED5);
//hidden: LED5
assign LED5 = IN;
endmodule
