module cOUT_PIN18(input wire OUT, output wire OUT_PIN18);
//hidden: OUT_PIN18
//position: 403,37,DE0nano
assign OUT_PIN18 = OUT;
endmodule
