module cLED3(input wire IN, output wire LED3);
//hidden: LED3
//position: 252,85,DE0nano
assign LED3 = IN;
endmodule
