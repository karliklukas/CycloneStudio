module cOUT_PIN11(input wire OUT, output wire OUT_PIN11);
//hidden: OUT_PIN11
//position: 129,302,DE0nano
assign OUT_PIN11 = OUT;
endmodule
