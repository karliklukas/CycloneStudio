module cOUT_PIN4(input wire OUT, output wire OUT_PIN4);
//hidden: OUT_PIN4
//position: 172,37,DE0nano;206,407,StormIV
assign OUT_PIN4 = OUT;
endmodule
