module cOUT_PIN19(input wire OUT, output wire OUT_PIN19);
//hidden: OUT_PIN19
//position: 403,51,DE0nano
assign OUT_PIN19 = OUT;
endmodule
