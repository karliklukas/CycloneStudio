module cKEY2(input wire KEY2, output wire OUT);
//hidden: KEY2
assign OUT = KEY2;
endmodule
