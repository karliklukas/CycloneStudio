module cOUT_PIN5(input wire OUT, output wire OUT_PIN5);
//hidden: OUT_PIN5
//position: 186,37,DE0nano;216,396,StormIV
assign OUT_PIN5 = OUT;
endmodule
