module cIN_PIN(input wire PIN, output wire IN);
//hidden: PIN
assign IN = PIN;
endmodule
