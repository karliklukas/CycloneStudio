module cIN_PIN16(input wire IN_PIN16, output wire IN);
//hidden: IN_PIN16
//position: 375,300,DE0nano
assign IN = IN_PIN16;
endmodule
