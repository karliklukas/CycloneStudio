module cvystup(input wire OUT, output wire vystup);
//hidden: vystup
assign vystup = OUT;
endmodule
