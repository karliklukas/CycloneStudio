module cOUT_PIN5(input wire OUT, output wire PIN5);
//hidden: PIN5
assign PIN5 = OUT;
endmodule
