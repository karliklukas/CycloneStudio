module cOUT_PIN9(input wire OUT, output wire OUT_PIN9);
//hidden: OUT_PIN9
assign OUT_PIN9 = OUT;
endmodule
