module cKEY_RESET(input wire KEY_RESET, output wire OUT);
//hidden: KEY_RESET
//position: 50,237,StormIV
assign OUT = KEY_RESET;
endmodule
