module cIN_PIN8(input wire PIN8, output wire IN);
//hidden: PIN8
assign IN = PIN8;
endmodule
