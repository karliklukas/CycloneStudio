module cLED3(input wire IN, output wire LED3);
//hidden: LED3
//position: 110,345,StormIV
assign LED3 = IN;
endmodule
