module cout1(input wire OUT, output wire out1);
//hidden: out1
assign out1 = OUT;
endmodule
