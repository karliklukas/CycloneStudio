module cOUT_vystup_a(input wire OUT, output wire vystup_a);
//hidden: vystup_a
assign vystup_a = OUT;
endmodule
