module cOUT_PIN8(input wire OUT, output wire OUT_PIN8);
//hidden: OUT_PIN8
assign OUT_PIN8 = OUT;
endmodule
