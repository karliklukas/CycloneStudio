module cLED0(input wire IN, output wire LED0);
//hidden: LED0
assign LED0 = IN;
endmodule
