module cLED7(input wire IN, output wire LED7);
//hidden: LED7
//position: 110,254,StormIV
assign LED7 = IN;
endmodule
