module cCLK_50MHz(input wire CLK_50MHz, output wire OUT);
//hidden: CLK_50MHz
assign OUT = CLK_50MHz;
endmodule
