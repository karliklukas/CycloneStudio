module cIN_PIN2(input wire IN_PIN2, output wire IN);
//hidden: IN_PIN2
//position: 144,300,DE0nano;259,196,StormIV
assign IN = IN_PIN2;
endmodule
