module cCustIn1(input wire CustIn1, output wire IN);
//hidden: CustIn1
assign IN = CustIn1;
endmodule
