module cLED3(input wire IN, output wire LED3);
//hidden: LED3
assign LED3 = IN;
endmodule
