module cOUT_PIN13(input wire OUT, output wire OUT_PIN13);
//hidden: OUT_PIN13
//position: 316,37,DE0nano
assign OUT_PIN13 = OUT;
endmodule
