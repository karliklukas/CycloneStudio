module cvystup_d(input wire OUT, output wire vystup_d);
//hidden: vystup_d
assign vystup_d = OUT;
endmodule
