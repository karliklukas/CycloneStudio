module cKEY1(input wire KEY1, output wire OUT);
//hidden: KEY1
//position: 340,89,DE0nano
assign OUT = KEY1;
endmodule
