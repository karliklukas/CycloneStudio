module cZERO(output wire Y);
assign Y = 1'b0;
endmodule
