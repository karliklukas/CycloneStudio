module cOUT_vystup_b(input wire OUT, output wire vystup_b);
//hidden: vystup_b
assign vystup_b = OUT;
endmodule
