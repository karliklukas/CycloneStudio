module cIN_PIN6(input wire PIN6, output wire IN);
//hidden: PIN6
assign IN = PIN6;
endmodule
