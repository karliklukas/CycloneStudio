module cIN_PIN10(input wire IN_PIN10, output wire IN);
//hidden: IN_PIN10
assign IN = IN_PIN10;
endmodule
