module cKEY2(input wire KEY2, output wire OUT);
//hidden: KEY2
//position: 50,367,StormIV
assign OUT = KEY2;
endmodule
