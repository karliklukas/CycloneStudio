module cIN_PIN3(input wire PIN3, output wire IN);
//hidden: PIN3
assign IN = PIN3;
endmodule
