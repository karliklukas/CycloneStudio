module cLED7(input wire IN, output wire LED7);
//hidden: LED7
//position: 183,85,DE0nano
assign LED7 = IN;
endmodule
