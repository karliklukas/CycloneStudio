module cIN_PIN7(input wire IN_PIN7, output wire IN);
//hidden: IN_PIN7
//position: 231,300,DE0nano;291,186,StormIV
assign IN = IN_PIN7;
endmodule
