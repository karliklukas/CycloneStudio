module cIN_PIN1(input wire IN_PIN1, output wire IN);
//hidden: IN_PIN1
//position: 129,300,DE0nano;259,186,StormIV
assign IN = IN_PIN1;
endmodule
