module cOUT_PIN12(input wire OUT, output wire OUT_PIN12);
//hidden: OUT_PIN12
//position: 302,37,DE0nano
assign OUT_PIN12 = OUT;
endmodule
