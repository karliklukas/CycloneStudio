module cIN_PIN18(input wire IN_PIN18, output wire IN);
//hidden: IN_PIN18
//position: 404,300,DE0nano
assign IN = IN_PIN18;
endmodule
