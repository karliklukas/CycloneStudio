module cpoiu(input wire poiu, output wire IN);
//hidden: poiu
assign IN = poiu;
endmodule
