module cOUT_PIN1(input wire OUT, output wire PIN1);
//hidden: PIN1
assign PIN1 = OUT;
endmodule
