module cIN_PIN9(input wire IN_PIN9, output wire IN);
//hidden: IN_PIN9
assign IN = IN_PIN9;
endmodule
