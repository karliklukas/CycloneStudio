module cLED2(input wire IN, output wire LED2);
//hidden: LED2
//position: 269,85,DE0nano
assign LED2 = IN;
endmodule
