module cLED6(input wire IN, output wire LED6);
//hidden: LED6
//position: 200,85,DE0nano
assign LED6 = IN;
endmodule
