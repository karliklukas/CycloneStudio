module cLED1(input wire IN, output wire LED1);
//hidden: LED1
//position: 110,391,StormIV
assign LED1 = IN;
endmodule
