module cOUT_PIN2(input wire OUT, output wire PIN2);
//hidden: PIN2
assign PIN2 = OUT;
endmodule
