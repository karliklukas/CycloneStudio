module cvstup_D(input wire vstup_D, output wire IN);
//hidden: vstup_D
assign IN = vstup_D;
endmodule
