module cOUT_PIN12(input wire OUT, output wire OUT_PIN12);
//hidden: OUT_PIN12
assign OUT_PIN12 = OUT;
endmodule
