module cvystup3(input wire OUT, output wire vystup3);
//hidden: vystup3
assign vystup3 = OUT;
endmodule
