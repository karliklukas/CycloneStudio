module cOUT_PIN3(input wire OUT, output wire OUT_PIN3);
//hidden: OUT_PIN3
assign OUT_PIN3 = OUT;
endmodule
