module cKEYreset(input wire KEYreset, output wire OUT);
//hidden: KEYreset
assign OUT = KEYreset;
endmodule
