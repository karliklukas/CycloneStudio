module cOUT_PIN16(input wire OUT, output wire OUT_PIN16);
//hidden: OUT_PIN16
//position: 375,37,DE0nano
assign OUT_PIN16 = OUT;
endmodule
