module cIN_PIN18(input wire IN_PIN18, output wire IN);
//hidden: IN_PIN18
assign IN = IN_PIN18;
endmodule
