module cvstup_A(input wire vstup_A, output wire IN);
//hidden: vstup_A
assign IN = vstup_A;
endmodule
