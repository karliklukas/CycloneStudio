module cOUT_PIN3(input wire OUT, output wire OUT_PIN3);
//hidden: OUT_PIN3
//position: 157,37,DE0nano;206,396,StormIV
assign OUT_PIN3 = OUT;
endmodule
