module cvstupA(input wire vstupA, output wire IN);
//hidden: vstupA
assign IN = vstupA;
endmodule
