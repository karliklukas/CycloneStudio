module cIN_PIN1(input wire IN_PIN1, output wire IN);
//hidden: IN_PIN1
//position: 139,263,DE0nano;139,263,StormIV
assign IN = IN_PIN1;
endmodule
