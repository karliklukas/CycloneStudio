module cvstup(input wire vstup, output wire IN);
//hidden: vstup
assign IN = vstup;
endmodule
