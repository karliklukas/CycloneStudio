module cOUT_PIN15(input wire OUT, output wire OUT_PIN15);
//hidden: OUT_PIN15
assign OUT_PIN15 = OUT;
endmodule
