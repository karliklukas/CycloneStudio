module cOUT_PIN13(input wire OUT, output wire OUT_PIN13);
//hidden: OUT_PIN13
assign OUT_PIN13 = OUT;
endmodule
