module cIN_PIN3(input wire IN_PIN3, output wire IN);
//hidden: IN_PIN3
//position: 158,300,DE0nano;270,186,StormIV
assign IN = IN_PIN3;
endmodule
