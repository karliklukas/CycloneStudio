module cIN_PIN14(input wire IN_PIN14, output wire IN);
//hidden: IN_PIN14
assign IN = IN_PIN14;
endmodule
