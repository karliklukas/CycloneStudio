module cIN_PIN5(input wire IN_PIN5, output wire IN);
//hidden: IN_PIN5
assign IN = IN_PIN5;
endmodule
