module cLED4(input wire IN, output wire LED4);
//hidden: LED4
assign LED4 = IN;
endmodule
