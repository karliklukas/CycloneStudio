module cCst1(input wire Cst1, output wire IN);
//hidden: Cst1
assign IN = Cst1;
endmodule
