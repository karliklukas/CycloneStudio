module cvystup6(input wire OUT, output wire vystup6);
//hidden: vystup6
assign vystup6 = OUT;
endmodule
