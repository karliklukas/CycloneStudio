module cOUT_PIN10(input wire OUT, output wire OUT_PIN10);
//hidden: OUT_PIN10
//position: 273,37,DE0nano;238,407,StormIV
assign OUT_PIN10 = OUT;
endmodule
