module cIN_PIN1(input wire PIN1, output wire IN);
//hidden: PIN1
assign IN = PIN1;
endmodule
