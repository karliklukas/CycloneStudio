module ckjhkj(input wire OUT, output wire kjhkj);
//hidden: kjhkj
assign kjhkj = OUT;
endmodule
