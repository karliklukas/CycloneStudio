module cLED1(input wire IN, output wire LED1);
//hidden: LED1
assign LED1 = IN;
endmodule
