module cLED7(input wire IN, output wire LED7);
//hidden: LED7
assign LED7 = IN;
endmodule
