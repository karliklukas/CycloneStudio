module cKEY4(input wire KEY4, output wire OUT);
//hidden: KEY4
//position: 50,286,StormIV
assign OUT = KEY4;
endmodule
