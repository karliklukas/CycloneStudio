module cIN_PIN19(input wire IN_PIN19, output wire IN);
//hidden: IN_PIN19
//position: 129,283,DE0nano
assign IN = IN_PIN19;
endmodule
