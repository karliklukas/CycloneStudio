module cOUT_PIN10(input wire OUT, output wire OUT_PIN10);
//hidden: OUT_PIN10
assign OUT_PIN10 = OUT;
endmodule
