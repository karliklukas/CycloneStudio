module cIN_PIN7(input wire PIN7, output wire IN);
//hidden: PIN7
assign IN = PIN7;
endmodule
