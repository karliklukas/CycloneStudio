module cIN_PIN7(input wire IN_PIN7, output wire IN);
//hidden: IN_PIN7
assign IN = IN_PIN7;
endmodule
