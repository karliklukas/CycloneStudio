module cIN_PIN1(input wire IN_PIN1, output wire IN);
//hidden: IN_PIN1
assign IN = IN_PIN1;
endmodule
