module cvstup3(input wire vstup3, output wire IN);
//hidden: vstup3
assign IN = vstup3;
endmodule
