module cLED2(input wire IN, output wire LED2);
//hidden: LED2
assign LED2 = IN;
endmodule
