module cOUT_PIN9(input wire OUT, output wire OUT_PIN9);
//hidden: OUT_PIN9
//position: 259,37,DE0nano;238,396,StormIV
assign OUT_PIN9 = OUT;
endmodule
