module cOUT_PIN6(input wire OUT, output wire OUT_PIN6);
//hidden: OUT_PIN6
//position: 215,37,DE0nano;216,407,StormIV
assign OUT_PIN6 = OUT;
endmodule
