module cLED4(input wire IN, output wire LED4);
//hidden: LED4
//position: 110,322,StormIV
assign LED4 = IN;
endmodule
