module cLED5(input wire IN, output wire LED5);
//hidden: LED5
//position: 110,300,StormIV
assign LED5 = IN;
endmodule
