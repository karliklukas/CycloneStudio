module cvystup_c(input wire OUT, output wire vystup_c);
//hidden: vystup_c
assign vystup_c = OUT;
endmodule
