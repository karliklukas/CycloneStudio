module cIN_PIN6(input wire IN_PIN6, output wire IN);
//hidden: IN_PIN6
assign IN = IN_PIN6;
endmodule
