module cOUT_PIN(input wire OUT, output wire PIN);
//hidden: PIN
assign PIN = OUT;
endmodule
