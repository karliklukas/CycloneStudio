module cIN_PIN20(input wire IN_PIN20, output wire IN);
//hidden: IN_PIN20
//position: 144,283,DE0nano
assign IN = IN_PIN20;
endmodule
