module cOUT_PIN18(input wire OUT, output wire OUT_PIN18);
//hidden: OUT_PIN18
assign OUT_PIN18 = OUT;
endmodule
