module cIN_PIN17(input wire IN_PIN17, output wire IN);
//hidden: IN_PIN17
//position: 389,300,DE0nano
assign IN = IN_PIN17;
endmodule
