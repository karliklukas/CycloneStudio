module cCustIN(input wire CustIN, output wire IN);
//hidden: CustIN
assign IN = CustIN;
endmodule
