module cIN_PIN20(input wire IN_PIN20, output wire IN);
//hidden: IN_PIN20
assign IN = IN_PIN20;
endmodule
