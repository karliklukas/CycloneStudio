module cvystup2(input wire OUT, output wire vystup2);
//hidden: vystup2
assign vystup2 = OUT;
endmodule
