module coutLED1(input wire OUT, output wire outLED1);
//hidden: outLED1
assign outLED1 = OUT;
endmodule
