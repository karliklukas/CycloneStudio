module cvystup4(input wire OUT, output wire vystup4);
//hidden: vystup4
assign vystup4 = OUT;
endmodule
