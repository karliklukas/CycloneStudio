module cvystup8(input wire OUT, output wire vystup8);
//hidden: vystup8
assign vystup8 = OUT;
endmodule
