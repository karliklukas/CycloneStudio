module cOUT_PIN7(input wire OUT, output wire PIN7);
//hidden: PIN7
assign PIN7 = OUT;
endmodule
