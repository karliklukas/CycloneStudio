module cIN_PIN9(input wire PIN9, output wire IN);
//hidden: PIN9
assign IN = PIN9;
endmodule
