module cIN_PIN2(input wire IN_PIN2, output wire IN);
//hidden: IN_PIN2
assign IN = IN_PIN2;
endmodule
