module cIN_PIN11(input wire IN_PIN11, output wire IN);
//hidden: IN_PIN11
//position: 288,300,DE0nano
assign IN = IN_PIN11;
endmodule
