module cinRESET(input wire inRESET, output wire IN);
//hidden: inRESET
assign IN = inRESET;
endmodule
