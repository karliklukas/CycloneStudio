module cLED8(input wire IN, output wire LED8);
//hidden: LED8
//position: 110,232,StormIV
assign LED8 = IN;
endmodule
