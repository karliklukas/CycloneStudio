module cOUT_PIN11(input wire OUT, output wire OUT_PIN11);
//hidden: OUT_PIN11
assign OUT_PIN11 = OUT;
endmodule
