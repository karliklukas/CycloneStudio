module cOUT_PIN3(input wire OUT, output wire PIN3);
//hidden: PIN3
assign PIN3 = OUT;
endmodule
