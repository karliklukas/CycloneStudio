module cIN_PIN8(input wire IN_PIN8, output wire IN);
//hidden: IN_PIN8
//position: 245,300,DE0nano;291,196,StormIV
assign IN = IN_PIN8;
endmodule
