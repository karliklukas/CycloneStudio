module cIN_PIN15(input wire IN_PIN15, output wire IN);
//hidden: IN_PIN15
assign IN = IN_PIN15;
endmodule
