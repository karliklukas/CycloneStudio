module cOUT_PIN7(input wire OUT, output wire OUT_PIN7);
//hidden: OUT_PIN7
//position: 230,37,DE0nano;227,396,StormIV
assign OUT_PIN7 = OUT;
endmodule
