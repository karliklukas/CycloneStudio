module cIN_PIN8(input wire IN_PIN8, output wire IN);
//hidden: IN_PIN8
assign IN = IN_PIN8;
endmodule
