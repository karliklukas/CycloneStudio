module cOUT_PIN2(input wire OUT, output wire OUT_PIN2);
//hidden: OUT_PIN2
assign OUT_PIN2 = OUT;
endmodule
