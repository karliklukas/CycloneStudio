module cLED5(input wire IN, output wire LED5);
//hidden: LED5
//position: 217,85,DE0nano
assign LED5 = IN;
endmodule
