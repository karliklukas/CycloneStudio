module cIN_PIN9(input wire IN_PIN9, output wire IN);
//hidden: IN_PIN9
//position: 259,300,DE0nano;302,186,StormIV
assign IN = IN_PIN9;
endmodule
