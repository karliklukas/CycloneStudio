module cIN_vstup_C(input wire vstup_C, output wire IN);
//hidden: vstup_C
assign IN = vstup_C;
endmodule
