module cOUT_PIN4(input wire OUT, output wire PIN4);
//hidden: PIN4
assign PIN4 = OUT;
endmodule
