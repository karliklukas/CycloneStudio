module cOUT_PIN11(input wire OUT, output wire OUT_PIN11);
//hidden: OUT_PIN11
//position: 288,37,DE0nano
assign OUT_PIN11 = OUT;
endmodule
