module cvystup_e(input wire OUT, output wire vystup_e);
//hidden: vystup_e
assign vystup_e = OUT;
endmodule
