module cIN_PIN4(input wire PIN4, output wire IN);
//hidden: PIN4
assign IN = PIN4;
endmodule
