module cLED1(input wire IN, output wire LED1);
//hidden: LED1
//position: 287,85,DE0nano
assign LED1 = IN;
endmodule
