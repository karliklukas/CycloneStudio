module cIN_PIN4(input wire IN_PIN4, output wire IN);
//hidden: IN_PIN4
//position: 173,300,DE0nano;270,196,StormIV
assign IN = IN_PIN4;
endmodule
