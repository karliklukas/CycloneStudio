module cvstupB(input wire vstupB, output wire IN);
//hidden: vstupB
assign IN = vstupB;
endmodule
