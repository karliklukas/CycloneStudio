module cOUT_PIN6(input wire OUT, output wire OUT_PIN6);
//hidden: OUT_PIN6
assign OUT_PIN6 = OUT;
endmodule
