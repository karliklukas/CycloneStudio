module cOUT_PIN8(input wire OUT, output wire PIN8);
//hidden: PIN8
assign PIN8 = OUT;
endmodule
