module cIN_vstup_B(input wire vstup_B, output wire IN);
//hidden: vstup_B
assign IN = vstup_B;
endmodule
