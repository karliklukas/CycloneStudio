module cBeeper(input wire OUT, output wire Beeper);
//hidden: Beeper
//position: 90,481,StormIV
assign Beeper = OUT;
endmodule
