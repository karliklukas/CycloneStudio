module cIN_PIN5(input wire IN_PIN5, output wire IN);
//hidden: IN_PIN5
//position: 187,300,DE0nano;281,186,StormIV
assign IN = IN_PIN5;
endmodule
