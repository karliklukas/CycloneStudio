module cKEY3(input wire KEY3, output wire OUT);
//hidden: KEY3
//position: 50,326,StormIV
assign OUT = KEY3;
endmodule
