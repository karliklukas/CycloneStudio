module cIN_PIN10(input wire IN_PIN10, output wire IN);
//hidden: IN_PIN10
//position: 273,300,DE0nano;302,196,StormIV
assign IN = IN_PIN10;
endmodule
