module cAdsd(input wire Adsd, output wire IN);
//hidden: Adsd
assign IN = Adsd;
endmodule
