module cOUT_vystup_f(input wire OUT, output wire vystup_f);
//hidden: vystup_f
assign vystup_f = OUT;
endmodule
