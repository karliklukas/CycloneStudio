module cKEY0(input wire KEY0, output wire OUT);
//hidden: KEY0
//position: 380,89,DE0nano
assign OUT = KEY0;
endmodule
