module cIN_PIN10(input wire PIN10, output wire IN);
//hidden: PIN10
assign IN = PIN10;
endmodule
