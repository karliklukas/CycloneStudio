module cBeeper(input wire OUT, output wire Beeper);
//hidden: Beeper
assign Beeper = OUT;
endmodule
