module cKEY_RESET(input wire KEY_RESET, output wire OUT);
//hidden: KEY_RESET
assign OUT = KEY_RESET;
endmodule
