module cKEY1(input wire KEY1, output wire OUT);
//hidden: KEY1
//position: 50,408,StormIV
assign OUT = KEY1;
endmodule
