module cIN_PIN15(input wire IN_PIN15, output wire IN);
//hidden: IN_PIN15
//position: 361,300,DE0nano
assign IN = IN_PIN15;
endmodule
