module cvystup7(input wire OUT, output wire vystup7);
//hidden: vystup7
assign vystup7 = OUT;
endmodule
