module cvystup_g(input wire OUT, output wire vystup_g);
//hidden: vystup_g
assign vystup_g = OUT;
endmodule
