module cKEY1(input wire KEY1, output wire OUT);
//hidden: KEY1
assign OUT = KEY1;
endmodule
