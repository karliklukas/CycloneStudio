module cKEY4(input wire KEY4, output wire OUT);
//hidden: KEY4
assign OUT = KEY4;
endmodule
