module cOUT_PIN4(input wire OUT, output wire OUT_PIN4);
//hidden: OUT_PIN4
assign OUT_PIN4 = OUT;
endmodule
